    Mac OS X            	   2   �      �                                      ATTR ��   �   �   X                  �   X  com.apple.quarantine q/0000;5072fd5e;Google\x20Chrome;29FBEC83-47A8-4DA4-8AF1-9E28668E33A3|com.google.Chrome 