grammar dfa ;

synthesized attribute pp :: String ;

nonterminal Root with pp ;


